`ifndef APB_SEQ_ITEM_SVH
`define APB_SEQ_ITEM_SVH



`endif // APB_SEQ_ITEM_SVH