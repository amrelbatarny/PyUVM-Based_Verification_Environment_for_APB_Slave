bind APB_Wrapper APB_SVA APB_SVA_inst (.*);