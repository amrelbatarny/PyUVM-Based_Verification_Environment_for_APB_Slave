module dpi_exports;
    
    import APB_seq_item_pkg::*;

    


endmodule