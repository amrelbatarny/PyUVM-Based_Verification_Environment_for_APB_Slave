/***********************************************************************
 * Author : Amr El Batarny
 * File   : SVA_bind.sv
 * Brief  : Bindings for SystemVerilog assertions into the APB design.
 **********************************************************************/

bind APB_Wrapper APB_SVA APB_SVA_inst (.*);